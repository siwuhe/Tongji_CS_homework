`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Testbench for the top module (CPU + Memories)
//////////////////////////////////////////////////////////////////////////////////

module top_tb;

    // 1. ���嶥��ģ��������ź� (��������Ϊ reg)
    reg clk_in;
    reg enable;
    reg reset;
    reg start;

    // 2. ���嶥��ģ�������ź� (��������Ϊ wire)
    wire [7:0] o_seg;
    wire [7:0] o_sel;
    wire [7:0] i_addr;
     wire [15:0] result_f1_tb;
     wire [15:0] result_f2_tb;
     wire [15:0] result_f3_tb;
     wire [15:0] instruction;
    // ʱ�Ӳ���
    localparam CLK_PERIOD = 10; // 10ns ���� (100MHz)

    // 3. ʵ��������ģ��
    top uut (
        .clk_in(clk_in),
        .enable(enable),
        .reset(reset),
        .start(start),
        .o_seg(o_seg),
        .o_sel(o_sel),
        .i_addr(i_addr),
        .result_f1(result_f1_tb),
        .result_f2(result_f2_tb),
        .result_f3(result_f3_tb),
        .instruction(instruction)
    );

    // 4. ʱ�������߼�
    initial begin
        clk_in = 0;
        // ѭ������ʱ���ź�
        forever #(CLK_PERIOD / 2) clk_in = ~clk_in; 
    end

    // 5. �������� (��ʼ������λ������)
    initial begin
        // ��ʼ�����������ź�
        enable = 1'b0;
        reset  = 1'b0;
        start  = 1'b0;

        // �ȴ�ʱ���ȶ�
        @(posedge clk_in);

        // --- 1. ������λ ---
        // ȷ�����мĴ����ʹ洢����ʼ��
        reset  = 1'b1;
        enable = 1'b1; // ���� CPU ���ڴ湤��

        // ���ָ�λ 5 ������
        repeat(5) @(posedge clk_in);

        // --- 2. ������λ ---
        reset = 1'b0;
        $display("System Reset complete. Starting CPU.");

        // --- 3. ������������ ---
        start = 1'b1;
        @(posedge clk_in);
        start = 1'b0; // ����������� 1 ������

        // --- 4. ���з��� ---
        // �����㹻����ʱ�䣬�� CPU �������ˤ�����㷨
        repeat(500000) @(posedge clk_in); 

        // --- 5. ������� ---
        $display("Simulation finished. Final results should be in registers R14 and R15.");
        $finish; 
    end

    // ��ѡ�����ε����������� Vivado �в鿴�ڲ��ź�
    initial begin
        $dumpfile("top.vcd");
        $dumpvars(0, top_tb); 
    end
    
endmodule