`timescale 1ns / 1ps

module dmem(
    input clk,     
    input ram_ena, 
    input wena,    
    input [9 : 0] addr,     // ���ģ���ַλ��� 7:0 (8λ) ��Ϊ 9:0 (10λ)
    input [31 : 0] data_in,  // ���ģ�����λ��� 15:0 (16λ) ��Ϊ 31:0 (32λ)
    output [31 : 0] data_out // ���ģ�����λ��� 15:0 (16λ) ��Ϊ 31:0 (32λ)
    );
    
    // 1024 x 32-bit �洢�� (2^10 = 1024)
    // �洢�������� 256 �� 16λ�� ������ 1024 �� 32λ��
    reg [31:0] data [1023:0]; 
    
    // ---- �ڴ��ʼ�� ----
    integer i;
    initial begin
        // ȫ����ʼ��Ϊ 0��������� xxxx��
        // ѭ����Χ�� 256 ������ 1024
        for (i = 0; i < 1024; i = i + 1)
            data[i] = 32'h0000_0000; // ���ģ���ʼ��ֵҲ��Ϊ 32λ

        // ����ѡ��������Ĳ��Գ����ʼ��һЩ���ݣ�
        // data[10'h000] = 32'h0000_0080; // ʾ������ַ 0 �洢 32λֵ 0x80
    end
    
    // �첽��ȡ
    // ���ģ���ȡ����Ϊ 32λ��δ����ʱ��� 32λ����̬
    assign data_out = ram_ena ? data[addr] : 32'hzzzz_zzzz;
    
    // ͬ��д��
    always @ (posedge clk)
    begin
        if (ram_ena && wena)
            data[addr] <= data_in;
    end
endmodule