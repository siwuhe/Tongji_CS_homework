module imem(
    input [9:0] addr,         // 8λ��ַ����Ӧ���256��ָ��
    output [31:0] instr       // 16λָ�����
    );

    // ʹ�� Xilinx IP �� dist_mem_gen
    dist_mem_gen_0 instr_mem(
        .a(addr),             // ��ַ����
        .spo(instr)           // �������
    );

endmodule