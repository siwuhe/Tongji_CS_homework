`timescale 1ns / 1ps

module dmem(
    input clk,     
    input ram_ena, 
    input wena,    
    input [7 : 0] addr,    
    input [15 : 0] data_in,
    output [15 : 0] data_out
    );
    
    // 256 x 16-bit �洢��
    reg [15:0] data [255:0]; 
    
    // ---- �ڴ��ʼ�� ----
    integer i;
    initial begin
        // ȫ����ʼ��Ϊ 0��������� xxxx��
        for (i = 0; i < 256; i = i + 1)
            data[i] = 16'h0000;

        // ����ѡ��������Ĳ��Գ����ʼ��һЩ���ݣ�
        // ���� DMEM[0] �� N��
        // data[8'h00] = 16'h0080;  
    end
    
    // �첽��ȡ
    assign data_out = ram_ena ? data[addr] : 16'hzzzz;
    
    // ͬ��д��
    always @ (posedge clk)
    begin
        if (ram_ena && wena)
            data[addr] <= data_in;
    end
endmodule
