module imem(
    input [7:0] addr,         // 8λ��ַ����Ӧ���256��ָ��
    output [15:0] instr       // 16λָ�����
    );

    // ʹ�� Xilinx IP �� dist_mem_gen
    dist_mem_gen_0 instr_mem(
        .a(addr),             // ��ַ����
        .spo(instr)           // �������
    );

endmodule
