`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Top Module for Nexys4DDR
//////////////////////////////////////////////////////////////////////////////////

module top(
    input  clk_in,     // ϵͳʱ��
    input  enable,     // BTNU   - CPU ��ʹ�ܣ����뱣�ְ��£�
    input  reset,      // BTNC   - ��λ����һ�¼��ɣ�
    input  start,      // BTND   - ���� CPU����һ�£�
    output [7:0] o_seg,
    output [7:0] o_sel
);

    // ======== CPU <-> IMEM / DMEM �ź� ========
    wire [15:0] instruction;
    wire [15:0] datain;
    wire [7:0]  i_addr;
    wire [7:0]  d_addr;
    wire wena;
    wire [15:0] dataout;

    // ======================================================
    //                  CLOCK DIVIDER
    // ======================================================
    reg [24:0] cnt = 0;

    always @(posedge clk_in or posedge reset)
        if (reset)
            cnt <= 0;
        else
            cnt <= cnt + 1'b1;

    // clk_cpu = clk_in / 8 �� 12.5MHz �� ��ˮ���㹻��
    wire clk_cpu = cnt[24];

    // ======================================================
    //                  7-SEG DISPLAY
    // ��ʾ PC �� 8 λ + ָ��� 8 λ
    // ======================================================
    wire [15:0] seg_data ={8'b0000_0000, instruction};

    seg7x16 seg7_inst(
        .clk(clk_in),
        .reset(reset),
        .cs(1'b1),
        .i_data(seg_data),
        .o_seg(o_seg),
        .o_sel(o_sel)
    );

    // ======================================================
    //                      CPU
    // ======================================================
    pcpu cpu_inst(
        .clk(clk_cpu),
        .enable(enable),     // �����ɰ������ƣ�����д��
        .reset(reset),
        .start(start),
        .instruction(instruction),
        .datain(datain),
        .i_addr(i_addr),
        .d_addr(d_addr),
        .wena(wena),
        .dataout(dataout),
        .result_f1(), .result_f2(), .result_f3()
    );

    // ======================================================
    //                      IMEM
    // ======================================================
    imem imem_inst(
        .addr(i_addr),
        .instr(instruction)
    );

    // ======================================================
    //                      DMEM
    // ======================================================
    dmem dmem_inst(
        .clk(clk_cpu),
        .ram_ena(enable),   // ����д�����ⲿ enable ����
        .wena(wena),
        .addr(d_addr),
        .data_in(dataout),
        .data_out(datain)
    );

endmodule
